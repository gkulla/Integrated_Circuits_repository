*** SPICE deck for cell inverter_sim{sch} from library EE4570_2
*** Created on Mon Sep 21, 2015 19:45:41
*** Last revised on Mon Sep 21, 2015 20:01:57
*** Written on Mon Sep 21, 2015 20:03:43 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT EE4570_2__inverter FROM CELL inverter{sch}
.SUBCKT EE4570_2__inverter In Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Out In gnd gnd NMOS L=0.4U W=0.8U
Mpmos-4@0 Out In vdd vdd PMOS L=0.4U W=1.6U
.ENDS EE4570_2__inverter

.global gnd vdd

*** TOP LEVEL CELL: inverter_sim{sch}
Xinverter@0 net@0 net@1 EE4570_2__inverter

* Spice Code nodes in cell cell 'inverter_sim{sch}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VIN In 0 PULSE(1.8 0 0 100p 100p 10n 20n)
.TRAN 0 50n
.include C:\Electric\C5_models.txt
.END
