*** SPICE deck for cell XOR_sim{sch} from library prova_library4_Nand_lay
*** Created on Thu Nov 12, 2015 22:15:05
*** Last revised on Sun Nov 22, 2015 20:57:04
*** Written on Sun Nov 22, 2015 20:57:09 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT prova_library4_Nand_lay__XOR FROM CELL XOR{sch}
.SUBCKT prova_library4_Nand_lay__XOR A AXORB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@66 A gnd gnd n L=0.4U W=1U
Mnmos-4@1 AXORB B net@66 net@66 n L=0.4U W=1U
Mnmos-4@2 AXORB net@134 net@6 net@6 n L=0.4U W=1U
Mnmos-4@3 net@6 net@125 gnd gnd n L=0.4U W=1U
Mnmos-4@4 net@134 A gnd gnd n L=0.4U W=1U
Mnmos-4@5 net@125 B gnd gnd n L=0.4U W=1U
Mpmos-4@0 AXORB net@134 net@19 net@19 p L=0.4U W=2U
Mpmos-4@1 net@19 B vdd vdd p L=0.4U W=2U
Mpmos-4@2 net@24 A vdd vdd p L=0.4U W=2U
Mpmos-4@3 AXORB net@125 net@24 net@24 p L=0.4U W=2U
Mpmos-4@5 net@134 A vdd vdd p L=0.4U W=2U
Mpmos-4@6 net@125 B vdd vdd p L=0.4U W=2U

* Spice Code nodes in cell cell 'XOR{sch}'
**.incude C:\Electric\MODEL_MOS.txt
**VDD VDD 0 DC 5
**VGND GND 0 DC 0
**VB B 0 DC 0
**VA A 0 DC 5
**.tran 0 40n
.ENDS prova_library4_Nand_lay__XOR

.global gnd vdd

*** TOP LEVEL CELL: XOR_sim{sch}
XXOR@0 A AXORB B prova_library4_Nand_lay__XOR

* Spice Code nodes in cell cell 'XOR_sim{sch}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 0
.tran 0 40n
.END
