*** SPICE deck for cell inverter_video_sim{sch} from library ProvaVideo1
*** Created on Wed Sep 23, 2015 10:21:59
*** Last revised on Wed Sep 23, 2015 10:35:15
*** Written on Wed Sep 23, 2015 10:35:24 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ProvaVideo1__inverter_video FROM CELL inverter_video{sch}
.SUBCKT ProvaVideo1__inverter_video In Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out In gnd gnd nmos L=0.4U W=2U
Mpmos@0 vdd In Out vdd pmos L=0.4U W=4U
.ENDS ProvaVideo1__inverter_video

.global gnd vdd

*** TOP LEVEL CELL: inverter_video_sim{sch}
Xinverter@0 net@0 net@1 ProvaVideo1__inverter_video

* Spice Code nodes in cell cell 'inverter_video_sim{sch}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
Vin in 0 DC 0
.include C:\Electric\C5_models.txt
.DC Vin 0 5 1mV
.END
