*** SPICE deck for cell six_transistor_SRAM{lay} from library prova_library2_IRSIM
*** Created on Thu Dec 03, 2015 13:30:19
*** Last revised on Thu Dec 03, 2015 14:12:01
*** Written on Thu Dec 03, 2015 14:17:19 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: six_transistor_SRAM{lay}
Mnmos@0 gnd net@15 net@2 gnd N L=0.4U W=1U AS=1.767P AD=3.9P PS=5.333U PD=9.8U
Mnmos@1 net@15 net@2 gnd gnd N L=0.4U W=1U AS=3.9P AD=1.867P PS=9.8U PD=5.467U
Mnmos@2 net@15 vdd In gnd N L=0.4U W=1U AS=1.4P AD=1.867P PS=4.8U PD=5.467U
Mnmos@3 Out vdd net@2 gnd N L=0.4U W=1U AS=1.767P AD=1.4P PS=5.333U PD=4.8U
Mpmos@0 vdd net@15 net@2 vdd P L=0.4U W=2U AS=1.767P AD=4.8P PS=5.333U PD=10.8U
Mpmos@1 net@15 net@2 vdd vdd P L=0.4U W=2U AS=4.8P AD=1.867P PS=10.8U PD=5.467U

* Spice Code nodes in cell cell 'six_transistor_SRAM{lay}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
Vin in 0 DC 1.8
.TRAN 0 50n
.include C:\Electric\MODEL_MOS.txt
.END
