*** SPICE deck for cell D_flipflop{sch} from library prova_library4_Nand_lay
*** Created on Mon Nov 30, 2015 20:02:32
*** Last revised on Mon Nov 30, 2015 22:41:35
*** Written on Mon Nov 30, 2015 22:43:24 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT prova_library4_Nand_lay__NAND_2 FROM CELL NAND_2{sch}
.SUBCKT prova_library4_Nand_lay__NAND_2 A AnandB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 AnandB A net@12 net@12 N L=0.4U W=0.8U
Mnmos-4@1 net@12 B gnd gnd N L=0.4U W=0.8U
Mpmos-4@0 AnandB B vdd vdd P L=0.4U W=1.6U
Mpmos-4@1 AnandB A vdd vdd P L=0.4U W=1.6U

* Spice Code nodes in cell cell 'NAND_2{sch}'
**.incude C:\Electric\MODEL_MOS.txt
**VDD VDD 0 DC 5
**VGND GND 0 DC 0
**VB B 0 DC 5
**VA A 0 DC 5
**.tran 0 40n
.ENDS prova_library4_Nand_lay__NAND_2

*** SUBCIRCUIT prova_library4_Nand_lay__inverter FROM CELL inverter{sch}
.SUBCKT prova_library4_Nand_lay__inverter In Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Out In gnd gnd n L=0.4U W=0.8U
Mpmos-4@0 Out In vdd vdd p L=0.4U W=1.6U
.ENDS prova_library4_Nand_lay__inverter

.global gnd vdd

*** TOP LEVEL CELL: D_flipflop{sch}
XNAND_2@0 D net@49 CK prova_library4_Nand_lay__NAND_2
XNAND_2@1 CK net@62 net@25 prova_library4_Nand_lay__NAND_2
XNAND_2@2 net@49 Q !Q prova_library4_Nand_lay__NAND_2
XNAND_2@3 Q !Q net@62 prova_library4_Nand_lay__NAND_2
Xinverter@0 D net@25 prova_library4_Nand_lay__inverter

* Spice Code nodes in cell cell 'D_flipflop{sch}'
**VDD VDD 0 DC 1.8
**VGND GND 0 DC 0
**VD D 0 DC PWL REPEAT FOREVER(0 0 0.99n 0 1n 1.8 1.99n 1.8 2n 0)ENDREPEAT
**VCK CK 0 DC PWL REPEAT FOREVER(0 0 0.499n 0 0.5n 1.8 0.99n 1.8 1n 0)ENDREPEAT
**.tran 0 20ns
**.include C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VD D 0 DC PWL (0 0 0.499n 0 0.5n 1.8 2.499n 1.8 2.5n 0 6.499n 0 6.5n 1.8 8.499n 1.8 8.5n 0)
VCK CK 0 DC PWL REPEAT FOREVER(0 0 0.99n 0 1n 1.8 1.99n 1.8 2n 0)ENDREPEAT
.tran 0 20ns
.include C:\Electric\MODEL_MOS.txt
.END
