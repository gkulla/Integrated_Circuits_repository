*** SPICE deck for cell nand_sim{sch} from library nand_gate
*** Created on Tue Nov 24, 2015 00:08:51
*** Last revised on Tue Nov 24, 2015 00:10:23
*** Written on Tue Nov 24, 2015 00:10:31 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT nand_gate__nand_gate FROM CELL nand_gate:nand_gate{sch}
.SUBCKT nand_gate__nand_gate A B F vdd
** GLOBAL 0
** GLOBAL vdd
Mnmos-4_0 net_88 B 0 0 N L=0.7U W=3.5U
Mnmos-4_1 F A net_88 net_88 N L=0.7U W=3.5U
Mpmos-4_0 vdd B F vdd P L=0.7U W=3.5U
Mpmos-4_1 vdd A F vdd P L=0.7U W=3.5U
.ENDS nand_gate__nand_gate

.global 0 vdd

*** TOP LEVEL CELL: nand_gate:nand_sim{sch}
Xnand_gat_0 A B F vdd nand_gate__nand_gate

* Spice Code nodes in cell cell 'nand_gate:nand_sim{sch}'
vdd vdd 0 DC 3.3
vgnd gnd 0 DC 0
vinA A 0 pwl(0 0 1ns 0 2ns 3.3 3ns 3.3)
vinB B 0 pwl(0 0 1ns 3.3 2ns 0 3ns 3.3)
.trans 0  3ns
.include C:\Users\Parmanand\Desktop\Electric\MOSmodel.txt
.END
