*** SPICE deck for cell inverter_video{sch} from library ProvaVideo
*** Created on Wed Sep 23, 2015 10:04:03
*** Last revised on Wed Sep 23, 2015 10:18:54
*** Written on Wed Sep 23, 2015 10:19:12 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inverter_video{sch}
Mnmos@0 Out In gnd gnd nmos L=0.4U W=2U
Mpmos@0 vdd In Out vdd pmos L=0.4U W=4U

* Spice Code nodes in cell cell 'inverter_video{sch}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
.include C:\Electric\C5_models.txt
.DC Vin 0 5 1mV
.END
