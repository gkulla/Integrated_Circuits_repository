*** SPICE deck for cell AND_sim{sch} from library prova_library4_Nand_lay
*** Created on Wed Dec 02, 2015 17:48:04
*** Last revised on Wed Dec 02, 2015 17:50:43
*** Written on Wed Dec 02, 2015 17:50:47 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT prova_library4_Nand_lay__AND FROM CELL AND{sch}
.SUBCKT prova_library4_Nand_lay__AND A AANDB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@5 A net@105 net@105 N L=0.4U W=1U
Mnmos-4@1 net@105 B gnd gnd N L=0.4U W=1U
Mnmos-4@3 AANDB net@5 gnd gnd n L=0.4U W=1U
Mpmos-4@0 net@5 B vdd vdd P L=0.4U W=2U
Mpmos-4@1 net@5 A vdd vdd P L=0.4U W=2U
Mpmos-4@2 AANDB net@5 vdd vdd p L=0.4U W=2U

* Spice Code nodes in cell cell 'AND{sch}'
**.incude C:\Electric\MODEL_MOS.txt
**VDD VDD 0 DC 5
**VGND GND 0 DC 0
**VB B 0 DC 0
**VA A 0 DC 5
**.tran 0 40n
.ENDS prova_library4_Nand_lay__AND

.global gnd vdd

*** TOP LEVEL CELL: AND_sim{sch}
XAND@0 A Out B prova_library4_Nand_lay__AND

* Spice Code nodes in cell cell 'AND_sim{sch}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 5
.tran 0 40n
.END
