*** SPICE deck for cell 3Input_OR_sim{sch} from library prova_library4_Nand_lay
*** Created on Thu Nov 12, 2015 23:01:31
*** Last revised on Sun Nov 22, 2015 21:05:20
*** Written on Sun Nov 22, 2015 21:05:23 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT prova_library4_Nand_lay__3Input_OR FROM CELL 3Input_OR{sch}
.SUBCKT prova_library4_Nand_lay__3Input_OR A AorBorC B C
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@0 A gnd gnd N L=0.4U W=1U
Mnmos-4@1 net@0 B gnd gnd N L=0.4U W=1U
Mnmos-4@2 net@0 C gnd gnd N L=0.4U W=1U
Mnmos-4@3 AorBorC net@0 gnd gnd n L=0.4U W=1U
Mpmos-4@0 net@0 C net@95 net@95 P L=0.4U W=2U
Mpmos-4@1 net@95 B net@90 net@90 P L=0.4U W=2U
Mpmos-4@2 net@90 A vdd vdd P L=0.4U W=2U
Mpmos-4@3 AorBorC net@0 vdd vdd p L=0.4U W=2U
.ENDS prova_library4_Nand_lay__3Input_OR

.global gnd vdd

*** TOP LEVEL CELL: 3Input_OR_sim{sch}
X_3Input_O@0 A AorBorC B C prova_library4_Nand_lay__3Input_OR

* Spice Code nodes in cell cell '3Input_OR_sim{sch}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 5
VC C 0 DC 5
.incude C:\Electric\MODEL_MOS.txt
.tran 0 40n
.END
