*** SPICE deck for cell XOR_TG{lay} from library Project2
*** Created on Fri Nov 13, 2015 18:43:41
*** Last revised on Fri Nov 13, 2015 19:05:12
*** Written on Fri Nov 13, 2015 19:05:16 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no power connection for P-transistor wells in cell 'Project2:XOR_TG{lay}'
*** WARNING: no ground connection for N-transistor wells in cell 'Project2:XOR_TG{lay}'

*** TOP LEVEL CELL: Project2:XOR_TG{lay}
Mnmos@0 notA B OUT gnd n L=0.4U W=1U AS=4.35P AD=4.45P PS=11.2U PD=11.4U
Mnmos@1 A_1 notB_1 OUT gnd n L=0.4U W=1U AS=4.35P AD=4.45P PS=11.2U PD=11.4U
Mpmos@0 notA notB OUT vdd p L=0.4U W=2U AS=4.35P AD=4.45P PS=11.2U PD=11.4U
Mpmos@1 A_1 B_1 OUT vdd p L=0.4U W=2U AS=4.35P AD=4.45P PS=11.2U PD=11.4U

* Spice Code nodes in cell cell 'Project2:XOR_TG{lay}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VnotA notA 0 DC 1.8
VB B 0 DC 1.8
VnotB notB 0 DC 1.8
VA_1 A_1 0 DC 0
VB_1 B_1 0 DC 1.8
VnotB_1 notB_1 0 DC 0
.TRAN 0 50n
.include C:\Electric\MODEL_MOS.txt
.END
