*** SPICE deck for cell XOR{lay} from library prova_library4_Nand_lay
*** Created on Fri Nov 13, 2015 12:58:03
*** Last revised on Sun Nov 15, 2015 10:36:39
*** Written on Sun Nov 15, 2015 10:36:42 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: XOR{lay}
Mnmos@0 net@303 net@151 AXORB gnd n L=0.4U W=1U AS=1.825P AD=1.3P PS=4.8U PD=4.6U
Mnmos@1 AXORB B net@299 gnd n L=0.4U W=1U AS=0.5P AD=1.825P PS=2U PD=4.8U
Mnmos@2 net@299 A gnd gnd n L=0.4U W=1U AS=6.1P AD=0.5P PS=14.2U PD=2U
Mnmos@3 gnd net@59 net@5 gnd n L=0.4U W=1U AS=1.4P AD=6.1P PS=4.8U PD=14.2U
Mnmos@4 net@59 B gnd gnd n L=0.4U W=1U AS=6.1P AD=2.3P PS=14.2U PD=6U
Mnmos@6 gnd A net@151 gnd n L=0.4U W=1U AS=2.4P AD=6.1P PS=6.2U PD=14.2U
Mpmos@0 AXORB net@151 net@308 vdd p L=0.4U W=2U AS=0.9P AD=1.825P PS=2.9U PD=4.8U
Mpmos@1 net@308 B vdd vdd p L=0.4U W=2U AS=7.15P AD=0.9P PS=15.45U PD=2.9U
Mpmos@2 vdd A net@311 vdd p L=0.4U W=2U AS=1.1P AD=7.15P PS=3.1U PD=15.45U
Mpmos@3 net@311 net@59 AXORB vdd p L=0.4U W=2U AS=1.825P AD=1.1P PS=4.8U PD=3.1U
Mpmos@4 net@59 B vdd vdd p L=0.4U W=2U AS=7.15P AD=2.3P PS=15.45U PD=6U
Mpmos@6 vdd A net@151 vdd p L=0.4U W=2U AS=2.4P AD=7.15P PS=6.2U PD=15.45U

* Spice Code nodes in cell cell 'XOR{lay}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 0
.tran 0 40n
.END
