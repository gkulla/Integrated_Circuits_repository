*** SPICE deck for cell 4_input_NAND{lay} from library prova_library4_Nand_lay
*** Created on Thu Dec 03, 2015 15:14:45
*** Last revised on Thu Dec 03, 2015 15:41:27
*** Written on Thu Dec 03, 2015 15:41:30 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: 4_input_NAND{lay}
Mnmos@0 Out A net@0 gnd n L=0.4U W=1U AS=0.45P AD=2.18P PS=2.1U PD=5.24U
Mnmos@1 net@0 B net@34 gnd n L=0.4U W=1U AS=0.43P AD=0.45P PS=1.9U PD=2.1U
Mnmos@2 net@34 C net@35 gnd n L=0.4U W=1U AS=0.44P AD=0.43P PS=2U PD=1.9U
Mnmos@3 net@35 D gnd gnd n L=0.4U W=1U AS=8.7P AD=0.44P PS=21.4U PD=2U
Mpmos@0 Out A vdd vdd p L=0.4U W=2U AS=4.55P AD=2.18P PS=9.65U PD=5.24U
Mpmos@1 vdd B Out vdd p L=0.4U W=2U AS=2.18P AD=4.55P PS=5.24U PD=9.65U
Mpmos@2 Out C vdd vdd p L=0.4U W=2U AS=4.55P AD=2.18P PS=9.65U PD=5.24U
Mpmos@3 vdd D Out vdd p L=0.4U W=2U AS=2.18P AD=4.55P PS=5.24U PD=9.65U

* Spice Code nodes in cell cell '4_input_NAND{lay}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 5
VA A 0 DC 0
VC C 0 DC 0
VD D 0 DC 0
.tran 0 40n
.END
