*** SPICE deck for cell complex_logic_function{sch} from library Project2
*** Created on Tue Oct 13, 2015 17:12:51
*** Last revised on Wed Oct 28, 2015 22:33:50
*** Written on Wed Oct 28, 2015 22:35:11 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: complex_logic_function{sch}
Mnmos-4@0 net@277 A gnd gnd n L=0.4U W=1U
Mnmos-4@1 net@218 B gnd gnd n L=0.4U W=1U
Mnmos-4@2 net@218 net@284 gnd gnd n L=0.4U W=1U
Mnmos-4@3 Out net@277 net@218 net@218 n L=0.4U W=1U
Mnmos-4@4 Out B net@218 net@218 n L=0.4U W=1U
Mnmos-4@5 Out C net@360 net@360 n L=0.4U W=1U
Mnmos-4@6 net@360 net@266 gnd gnd n L=0.4U W=1U
Mnmos-4@7 net@266 D gnd gnd n L=0.4U W=1U
Mnmos-4@8 net@284 C gnd gnd n L=0.4U W=1U
Mpmos-4@9 net@277 A vdd vdd p L=0.4U W=2U
Mpmos-4@10 Out C net@252 net@252 p L=0.4U W=2U
Mpmos-4@11 Out net@266 net@252 net@252 p L=0.4U W=2U
Mpmos-4@12 net@252 B net@412 net@412 p L=0.4U W=2U
Mpmos-4@13 net@412 net@277 vdd vdd p L=0.4U W=2U
Mpmos-4@14 net@432 B vdd vdd p L=0.4U W=2U
Mpmos-4@15 net@252 net@284 net@432 net@432 p L=0.4U W=2U
Mpmos-4@16 net@266 D vdd vdd p L=0.4U W=2U
Mpmos-4@17 net@284 C vdd vdd p L=0.4U W=2U

* Spice Code nodes in cell cell 'complex_logic_function{sch}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VA A 0 DC 1.8
VB B 0 DC 0
VD D 0 DC 0
VC C 0 Pulse(1.8 0 0 20n 40n 0.5u 1u)
**VD D 0 DC 0
.tran 0 3u
.include C:\Electric\MODEL_MOS.txt
.END
