*** SPICE deck for cell inverter_videos{ic} from library ProvaVideo
*** Created on Wed Sep 23, 2015 10:45:37
*** Last revised on Wed Sep 23, 2015 12:03:18
*** Written on Wed Sep 23, 2015 12:03:34 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: inverter_videos{ic}

* Spice Code nodes in cell cell 'inverter_videos{ic}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
Vin in 0 DC 0
.include C:\Electric\C5_models.txt
.DC Vin 0 5 1mV
.END
