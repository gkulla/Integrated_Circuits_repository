*** SPICE deck for cell D_vs_VBS_PMOS{sch} from library prova_library4_Nand_lay
*** Created on Tue Nov 03, 2015 19:21:06
*** Last revised on Tue Nov 03, 2015 19:38:24
*** Written on Wed Nov 04, 2015 20:25:37 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd
*** WARNING: no power connection for P-transistor wells in cell 'D_vs_VBS_PMOS{sch}'

*** TOP LEVEL CELL: D_vs_VBS_PMOS{sch}
Mpmos-4@0 net@5 net@0 gnd net@3 p L=0.4U W=2U
VVBS net@3 gnd DC 0V
VVSD gnd net@5 DC 2V
VVSG gnd net@0 DC 0V

* Spice Code nodes in cell cell 'D_vs_VBS_PMOS{sch}'
VGND GND 0 DC 0
.dc VVSG 0 5 1m VVBS 0 5 1
.incude C:\Electric\MODEL_MOS.txt
.END
