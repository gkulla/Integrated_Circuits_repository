*** SPICE deck for cell inverter_videos_sim{sch} from library ProvaVideo2
*** Created on Wed Sep 23, 2015 12:05:21
*** Last revised on Wed Sep 23, 2015 12:20:00
*** Written on Wed Sep 23, 2015 12:20:10 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ProvaVideo2__inverter_videos FROM CELL inverter_videos{sch}
.SUBCKT ProvaVideo2__inverter_videos In Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out In gnd gnd nmos L=0.4U W=2U
Mpmos@0 vdd In Out vdd pmos L=0.4U W=4U
.ENDS ProvaVideo2__inverter_videos

.global gnd vdd

*** TOP LEVEL CELL: inverter_videos_sim{sch}
Xinverter@0 In Out ProvaVideo2__inverter_videos

* Spice Code nodes in cell cell 'inverter_videos_sim{sch}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
Vin in 0 DC 0
.include C:\Electric\C5_models.txt
.DC Vin 0 5 1mV
.END
