*** SPICE deck for cell Dynamic4InputNand{lay} from library prova_library4_Nand_lay
*** Created on Sun Nov 08, 2015 16:56:29
*** Last revised on Sun Nov 08, 2015 17:25:31
*** Written on Sun Nov 08, 2015 17:25:40 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: Dynamic4InputNand{lay}
Mnmos@0 net@1 In1 Out gnd n L=0.4U W=1U AS=2.25P AD=0.43P PS=6U PD=1.9U
Mnmos@1 net@0 In2 net@1 gnd n L=0.4U W=1U AS=0.43P AD=0.43P PS=1.9U PD=1.9U
Mnmos@2 net@2 In3 net@0 gnd n L=0.4U W=1U AS=0.43P AD=0.45P PS=1.9U PD=1.9U
Mnmos@3 net@3 In4 net@2 gnd n L=0.4U W=1U AS=0.45P AD=0.44P PS=1.9U PD=2U
Mnmos@4 gnd CLK net@3 gnd n L=0.4U W=1U AS=0.44P AD=3.6P PS=2U PD=11.2U
Mpmos@0 vdd CLK Out vdd p L=0.4U W=2U AS=2.25P AD=7.4P PS=6U PD=17.8U

* Spice Code nodes in cell cell 'Dynamic4InputNand{lay}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VIn1 In1 0 DC 1.8
VIn2 In2 0 DC 1.8
VIn3 In3 0 DC 1.8
VIn4 In4 0 DC 1.8
VCLK CLK 0 Pulse(1.8 0 0 100p 100p 10n 20n)
.incude C:\Electric\MODEL_MOS.txt
.tran 0 50n
.END
