*** SPICE deck for cell inverter_serie{sch} from library prova_library2_IRSIM
*** Created on Wed Oct 14, 2015 23:27:12
*** Last revised on Thu Oct 15, 2015 15:23:27
*** Written on Thu Oct 15, 2015 15:23:32 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: prova_library2_IRSIM:inverter_serie{sch}
Mnmos-4@0 net@24 In gnd gnd n L=0.4U W=0.8U
Mnmos-4@1 Out net@24 gnd gnd n L=0.4U W=0.8U
Mpmos-4@0 net@24 In vdd vdd p L=0.4U W=0.8U
Mpmos-4@1 Out net@24 vdd vdd p L=0.4U W=0.8U

* Spice Code nodes in cell cell 'prova_library2_IRSIM:inverter_serie{sch}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
Vin in 0 Pulse(1.8 0 0 100p 100p 10n 20n)
**cload Out 0 1025fF
.TRAN 0 50n
.include C:\Electric\MODEL_MOS.txt
.END
