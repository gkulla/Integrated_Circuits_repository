*** SPICE deck for cell NAND_2{sch} from library prova_library4_Nand_lay
*** Created on Sun Sep 27, 2015 16:40:20
*** Last revised on Tue Nov 24, 2015 21:06:17
*** Written on Tue Nov 24, 2015 21:06:22 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: NAND_2{sch}
Mnmos-4@0 AnandB A net@12 net@12 N L=0.4U W=0.8U
Mnmos-4@1 net@12 B gnd gnd N L=0.4U W=0.8U
Mpmos-4@0 AnandB B vdd vdd P L=0.4U W=1.6U
Mpmos-4@1 AnandB A vdd vdd P L=0.4U W=1.6U

* Spice Code nodes in cell cell 'NAND_2{sch}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 5
VA A 0 DC 5
.tran 0 40n
.END
