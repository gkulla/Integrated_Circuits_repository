*** SPICE deck for cell Or_7inputs{sch} from library prova_library4_Nand_lay
*** Created on Sun Dec 13, 2015 18:08:37
*** Last revised on Sun Dec 13, 2015 18:15:02
*** Written on Sun Dec 13, 2015 18:15:07 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Or_7inputs{sch}
Mnmos-4@0 net@1 E gnd gnd N L=0.7U W=1.75U
Mnmos-4@1 net@1 F gnd gnd N L=0.7U W=1.75U
Mnmos-4@2 Out net@1 gnd gnd n L=0.7U W=1.75U
Mnmos-4@3 net@1 D gnd gnd N L=0.7U W=1.75U
Mnmos-4@4 net@1 C gnd gnd N L=0.7U W=1.75U
Mnmos-4@5 net@1 B gnd gnd N L=0.7U W=1.75U
Mnmos-4@6 net@1 A gnd gnd N L=0.7U W=1.75U
Mnmos-4@7 net@1 G gnd gnd N L=0.7U W=1.75U
Mpmos-4@0 net@6 D net@53 net@53 P L=0.7U W=3.5U
Mpmos-4@1 net@53 C net@29 net@29 P L=0.7U W=3.5U
Mpmos-4@2 net@29 B net@2 net@2 P L=0.7U W=3.5U
Mpmos-4@3 Out net@1 vdd vdd p L=0.7U W=3.5U
Mpmos-4@4 net@30 E net@6 net@6 P L=0.7U W=3.5U
Mpmos-4@5 net@132 F net@30 net@30 P L=0.7U W=3.5U
Mpmos-4@6 net@2 A vdd vdd P L=0.7U W=3.5U
Mpmos-4@8 net@1 G net@132 net@132 P L=0.7U W=3.5U

* Spice Code nodes in cell cell 'Or_7inputs{sch}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 0
VC C 0 DC 0
VD D 0 DC 0
VE E 0 DC 0
VF F 0 DC 0
.incude C:\Electric\MODEL_MOS.txt
.tran 0 40n
.END
