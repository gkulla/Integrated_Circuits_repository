*** SPICE deck for cell 6input_andgate{sch} from library 4input_andgate
*** Created on Sun Dec 13, 2015 21:43:13
*** Last revised on Mon Dec 14, 2015 09:37:01
*** Written on Mon Dec 14, 2015 10:28:03 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 4input_andgate:6input_andgate{sch}
Mnmos@0 net@49 D net@41 gnd N L=0.7U W=1.75U
Mnmos@1 net@36 C net@49 gnd N L=0.7U W=1.75U
Mnmos@2 net@3 B net@36 gnd N L=0.7U W=1.75U
Mnmos@3 net@0 A net@3 gnd N L=0.7U W=1.75U
Mnmos@4 Out net@0 gnd gnd N L=0.7U W=1.75U
Mnmos@5 net@41 E net@68 gnd N L=0.7U W=1.75U
Mnmos@6 net@68 F gnd gnd N L=0.7U W=1.75U
Mpmos@0 vdd A net@0 vdd P L=0.7U W=3.5U
Mpmos@1 vdd B net@0 vdd P L=0.7U W=3.5U
Mpmos@2 vdd C net@0 vdd P L=0.7U W=3.5U
Mpmos@3 vdd D net@0 vdd P L=0.7U W=3.5U
Mpmos@4 vdd net@0 Out vdd P L=0.7U W=3.5U
Mpmos@5 vdd E net@0 vdd P L=0.7U W=3.5U
Mpmos@6 vdd F net@0 vdd P L=0.7U W=3.5U

* Spice Code nodes in cell cell '4input_andgate:6input_andgate{sch}'
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VC C 0 DC 5
VB B 0 DC 5
VA A 0 DC 5
VD D 0 DC 5
VE E 0 DC 5
VF F 0 DC 5
.tran 0 40n
.END
