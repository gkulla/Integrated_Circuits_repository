*** SPICE deck for cell hwsix_cas{sch} from library prova_library2_IRSIM
*** Created on Mon Nov 30, 2015 18:34:48
*** Last revised on Mon Nov 30, 2015 19:10:51
*** Written on Mon Nov 30, 2015 19:12:27 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: hwsix_cas{sch}
Mnmos-4@1 net@51 A net@18 net@18 n L=0.4U W=1U
Mnmos-4@3 net@18 B net@9 net@9 n L=0.4U W=1U
Mnmos-4@5 net@9 CK gnd gnd n L=0.4U W=1U
Mnmos-4@6 net@47 net@51 gnd gnd n L=0.4U W=1U
Mnmos-4@7 net@97 net@47 net@81 net@81 n L=0.4U W=1U
Mnmos-4@8 net@97 C net@91 net@91 n L=0.4U W=1U
Mnmos-4@10 net@91 D net@81 net@81 n L=0.4U W=1U
Mnmos-4@11 net@81 CK gnd gnd n L=0.4U W=1U
Mnmos-4@12 Out net@97 gnd gnd n L=0.4U W=1U
Mpmos-4@0 net@51 CK vdd vdd n L=0.4U W=2U
Mpmos-4@2 net@47 net@51 vdd vdd n L=0.4U W=2U
Mpmos-4@3 net@97 CK vdd vdd n L=0.4U W=2U
Mpmos-4@4 Out net@97 vdd vdd n L=0.4U W=2U

* Spice Code nodes in cell cell 'hwsix_cas{sch}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VA A 0 DC PWL REPEAT FOREVER(0 0 7.99n 0 8n 1.8 15.99n 1.8 16n 0)ENDREPEAT
VB B 0 DC PWL REPEAT FOREVER(0 0 3.99n 0 4n 1.8 7.99n 1.8 8n 0)ENDREPEAT
VC C 0 DC PWL REPEAT FOREVER(0 0 1.99n 0 2n 1.8 3.99n 1.8 4n 0)ENDREPEAT
VD D 0 DC PWL REPEAT FOREVER(0 0 0.99n 0 1n 1.8 1.99n 1.8 2n 0)ENDREPEAT
VCK CK 0 DC PWL REPEAT FOREVER(0 0 0.499n 0 0.5n 1.8 0.7499n 1.8 0.75n 0)ENDREPEAT
.tran 0 20ns
.include C:\Electric\MODEL_MOS.txt
.END
