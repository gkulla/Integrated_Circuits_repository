*** SPICE deck for cell inverter_sim{sch} from library Indipendent_Study
*** Created on Fri Jul 21, 2017 21:13:18
*** Last revised on Thu Jul 27, 2017 11:10:04
*** Written on Thu Jul 27, 2017 11:10:11 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Indipendent_Study__inverter FROM CELL inverter{sch}
.SUBCKT Indipendent_Study__inverter in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=6U
.ENDS Indipendent_Study__inverter

.global gnd vdd

*** TOP LEVEL CELL: inverter_sim{sch}
Xinverter@0 in out Indipendent_Study__inverter

* Spice Code nodes in cell cell 'inverter_sim{sch}'
vdd vdd 0 DC 5
VGND GND 0 DC 0
vin in 0 PULSE(5 0 0 100p 100p 10n 20n)
.tran 0 50n
.include C:\Electric\panic\C5_models.txt
.END
