*** SPICE deck for cell Inv_20_10{sch} from library CMOSedu_1
*** Created on Sat Sep 05, 2015 15:29:06
*** Last revised on Sun Sep 06, 2015 14:58:25
*** Written on Mon Sep 07, 2015 11:46:11 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Inv_20_10{sch}
Mnmos@0 OUT IN gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd IN OUT vdd PMOS L=0.4U W=4U
Vin IN gnd DC 0V

* Spice Code nodes in cell cell 'Inv_20_10{sch}'
VDD VDD 0 DC 5
Vgnd GND 0 DC 0
.include C:\Electric\C5_models.txt
.DC Vin 0 5 1mV
.END
