*** SPICE deck for cell NOR{ic} from library prova_library4_Nand_lay
*** Created on Tue Nov 03, 2015 17:24:58
*** Last revised on Wed Dec 02, 2015 17:45:25
*** Written on Wed Dec 02, 2015 17:45:32 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NOR{ic}

* Spice Code nodes in cell cell 'NOR{ic}'
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 5
VA A 0 DC 0
.incude C:\Electric\MODEL_MOS.txt
.tran 0 40n
.END
