*** SPICE deck for cell AND{sch} from library prova_library4_Nand_lay
*** Created on Thu Nov 12, 2015 22:21:39
*** Last revised on Wed Dec 02, 2015 22:30:43
*** Written on Wed Dec 02, 2015 22:34:41 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: AND{sch}
Mnmos@0 net@128 B gnd gnd n L=0.4U W=1U
Mnmos@1 net@21 A net@128 gnd n L=0.4U W=1U
Mnmos@2 AANDB net@21 gnd gnd n L=0.4U W=1U
Mpmos@0 vdd net@21 AANDB vdd p L=0.4U W=2U
Mpmos@1 vdd A net@21 vdd p L=0.4U W=2U
Mpmos@2 vdd B net@21 vdd p L=0.4U W=2U

* Spice Code nodes in cell cell 'AND{sch}'
**.incude C:\Electric\MODEL_MOS.txt
**VDD VDD 0 DC 5
**VGND GND 0 DC 0
**VB B 0 DC 0
**VA A 0 DC 5
**.tran 0 40n
.incude C:\Electric\MODEL_MOS.txt
VDD VDD 0 DC 5
VGND GND 0 DC 0
VB B 0 DC 0
VA A 0 DC 5
.tran 0 40n
.END
