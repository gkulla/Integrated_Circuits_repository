*** SPICE deck for cell hwsix_cascade{sch} from library prova_library2_IRSIM
*** Created on Mon Nov 30, 2015 21:09:31
*** Last revised on Mon Nov 30, 2015 21:17:58
*** Written on Mon Nov 30, 2015 21:18:54 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: hwsix_cascade{sch}
Mnmos-4@0 net@42 A net@71 net@71 n L=0.4U W=1U
Mnmos-4@2 net@71 B net@22 net@22 n L=0.4U W=1U
Mnmos-4@4 net@22 CK gnd gnd n L=0.4U W=1U
Mnmos-4@5 net@29 net@42 gnd gnd n L=0.4U W=1U
Mnmos-4@6 net@83 net@29 net@99 net@99 n L=0.4U W=1U
Mnmos-4@7 net@83 C net@126 net@126 n L=0.4U W=1U
Mnmos-4@9 net@126 D net@99 net@99 n L=0.4U W=1U
Mnmos-4@10 net@99 net@96 gnd gnd n L=0.4U W=1U
Mnmos-4@11 Out net@83 gnd gnd n L=0.4U W=1U
Mpmos-4@0 net@42 CK vdd vdd n L=0.4U W=2U
Mpmos-4@2 net@29 net@42 vdd vdd n L=0.4U W=2U
Mpmos-4@3 net@83 net@96 vdd vdd n L=0.4U W=2U
Mpmos-4@4 Out net@83 vdd vdd n L=0.4U W=2U

* Spice Code nodes in cell cell 'hwsix_cascade{sch}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VA A 0 DC PWL REPEAT FOREVER(0 0 7.99n 0 8n 1.8 15.99n 1.8 16n 0)ENDREPEAT
VB B 0 DC PWL REPEAT FOREVER(0 0 3.99n 0 4n 1.8 7.99n 1.8 8n 0)ENDREPEAT
VC C 0 DC PWL REPEAT FOREVER(0 0 1.99n 0 2n 1.8 3.99n 1.8 4n 0)ENDREPEAT
VD D 0 DC PWL REPEAT FOREVER(0 0 0.99n 0 1n 1.8 1.99n 1.8 2n 0)ENDREPEAT
VCK CK 0 DC PWL REPEAT FOREVER(0 0 0.499n 0 0.5n 1.8 0.99n 1.8 1n 0)ENDREPEAT
.tran 0 20ns
.include C:\Electric\MODEL_MOS.txt
.END
