*** SPICE deck for cell hwsix{lay} from library prova_library2_IRSIM
*** Created on Mon Nov 30, 2015 20:56:29
*** Last revised on Wed Dec 02, 2015 21:25:21
*** Written on Wed Dec 02, 2015 21:25:25 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: hwsix{lay}
Mnmos@0 net@43 C Out gnd n L=0.4U W=1U AS=1.633P AD=0.5P PS=4.267U PD=2U
Mnmos@1 Out A net@11 gnd n L=0.4U W=1U AS=0.45P AD=1.633P PS=1.9U PD=4.267U
Mnmos@2 gnd CK net@0 gnd n L=0.4U W=1U AS=1P AD=3.2P PS=3U PD=10.4U
Mnmos@3 net@11 B net@10 gnd n L=0.4U W=1U AS=1.5P AD=0.45P PS=5U PD=1.9U
Mnmos@4 net@0 D net@43 gnd n L=0.4U W=1U AS=0.5P AD=1P PS=2U PD=3U
Mpmos@0 Out CK vdd vdd p L=0.4U W=2U AS=7.4P AD=1.633P PS=17.8U PD=4.267U

* Spice Code nodes in cell cell 'hwsix{lay}'
VDD VDD 0 DC 1.8
VGND GND 0 DC 0
VA A 0 DC PWL REPEAT FOREVER(0 0 15.99n 0 16n 1.8 31.99n 1.8 32n 0)ENDREPEAT
VB B 0 DC PWL REPEAT FOREVER(0 0 7.99n 0 8n 1.8 15.99n 1.8 16n 0)ENDREPEAT
VC C 0 DC PWL REPEAT FOREVER(0 0 3.99n 0 4n 1.8 7.99n 1.8 8n 0)ENDREPEAT
VD D 0 DC PWL REPEAT FOREVER(0 0 1.99n 0 2n 1.8 3.99n 1.8 4n 0)ENDREPEAT
VCK CK 0 DC PWL REPEAT FOREVER(0 0 0.99n 0 1n 1.8 1.99n 1.8 2n 0)ENDREPEAT
.tran 0 70ns
.include C:\Electric\MODEL_MOS.txt
.END
